RC Low-Pass Filter
* Simple 1st-order RC low-pass, f_3dB ≈ 15.9 kHz
Vin in 0 AC 1
R1 in out 1k
C1 out 0 10n
.ac dec 50 1 100MEG
.meas ac f3dB WHEN vdb(out)=-3 FALL=1
.end
