RC Low-Pass — R Sweep
* Demonstrates .step param sweep: R from 500 to 2k in 500 steps
Vin in 0 AC 1
R1 in out {Rval}
C1 out 0 10n
.param Rval=1k
.step param Rval 500 2000 500
.ac dec 50 1 100MEG
.meas ac f3dB WHEN vdb(out)=-3 FALL=1
.end
